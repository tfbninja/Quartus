module mux7(input [6:0] x, input [6:0] off, input enable);
	
endmodule
