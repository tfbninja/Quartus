module L4_P3(

	//////////// LED //////////
	output [1:0]LEDR,

	//////////// SW //////////
	input [9:0]SW
);



//=======================================================
//  REG/WIRE declarations
//=======================================================
	wire [1:0]a, [1:0]b, [1:0]c, x, y;
	assign x = SW[9];
	assign y = SW[8];
	

//=======================================================
//  Structural coding
//=======================================================
	assign LEDR[9] = x;
	assign LEDR[8] = y;
	assign LEDR[1:0] = 

endmodule
